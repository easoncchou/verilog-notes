`include "fifo_mem.v"
// timescale directive: time unit / time precision for simulations
`timescale 10 ps / 10 ps
// preprocessor directive
`define DELAY 10 // define micro with value 10 as a parameter

module tb_fifo_32;

// parameter definitions
parameter ENDTIME = 40000;

// DUT Input Regs

// DUT Output Wires

// DUT Instantiation

// Initial Conditions

// Generating Test Vectors

// Debug FIFO

// Self-Checking

// Determine the simulation limit

endmodule